
module vini

